interface (clk,rst);
endinterface
